/*
`timescale 1ns/1ps
`include "UART_TX.v"
`include "UART_RX.v"
`include "LFSR.v"
`include "SAR.v"

module UART_TB;

  // Clock and reset
  reg r_Clock = 0;
  reg r_Rst_L = 1;

  // UART signals
  reg r_TX_DV = 0;
  wire [7:0] w_LFSR_Byte;
  wire w_TX_Serial;
  wire w_RX_DV;
  wire [7:0] w_RX_Byte;
  wire [15:0] w_SAR_Tx;
  wire [15:0] w_SAR_Rx;

  // Instantiate the UART modules
  UART_TX #(.CLK_FREQ(25000000), .BAUD_RATE(115200)) UART_TX_INST (
    .i_Rst_L(r_Rst_L),
    .i_Clock(r_Clock),
    .i_TX_DV(r_TX_DV),
    .i_TX_Byte(w_LFSR_Byte),
    .o_TX_Active(),
    .o_TX_Serial(w_TX_Serial),
    .o_TX_Done()
  );

  UART_RX #(.CLK_FREQ(25000000), .BAUD_RATE(115200)) UART_RX_INST (
    .i_Clock(r_Clock),
    .i_RX_Serial(w_TX_Serial),
    .o_RX_DV(w_RX_DV),
    .o_RX_Byte(w_RX_Byte)
  );

  LFSR #(.WIDTH(16), .SEED(16'hACE1)) LFSR_INST (
    .i_Clock(r_Clock),
    .i_Enable(r_TX_DV),
    .o_LFSR_Byte(w_LFSR_Byte)
  );

  SAR #(.WIDTH(16)) SAR_TX_INST (
    .i_Clock(r_Clock),
    .i_Enable(r_TX_DV),
    .i_Data(w_LFSR_Byte),
    .o_SAR(w_SAR_Tx)
  );

  SAR #(.WIDTH(16)) SAR_RX_INST (
    .i_Clock(r_Clock),
    .i_Enable(w_RX_DV),
    .i_Data(w_RX_Byte),
    .o_SAR(w_SAR_Rx)
  );

  // Clock generation
  always #10 r_Clock = ~r_Clock;  // 50MHz clock
    integer i;
  // Main Testing:
  initial
  begin


    // Open a VCD file for waveform analysis
    $dumpfile("dump.vcd");
    $dumpvars(0, UART_TB);
    $dumpvars(1, UART_TX_INST);
    $dumpvars(1, UART_RX_INST);

    // Apply reset
    r_Rst_L = 1'b0;
    #100;
    r_Rst_L = 1'b1;
    #100;

    for (i = 0; i < 10; i = i + 1) begin
      $display("Starting iteration %0d", i);
      // Tell UART to send a command (exercise TX)
      @(posedge r_Clock);
      @(posedge r_Clock);
      r_TX_DV   <= 1'b1;
      @(posedge r_Clock);
      r_TX_DV <= 1'b0;

      // Wait for the data to be received
      wait (w_RX_DV);

      // Debug: print values for each iteration
      $display("LFSR Byte Sent: %h", w_LFSR_Byte);
      $display("Received Byte: %h", w_RX_Byte);

      // Check that the correct command was received
      if (w_RX_Byte !== w_LFSR_Byte)
        $display("Test Failed - Incorrect Byte Received. Expected: %h, Received: %h", w_LFSR_Byte, w_RX_Byte);
      else
        $display("Test Passed - Correct Byte Received. Byte: %h", w_RX_Byte);
        
      #100000; // Add delay between iterations to ensure proper timing
    end

    // Check final SAR values
    if (w_SAR_Tx === w_SAR_Rx)
      $display("Test Passed - Signatures Match. SAR_Tx: %h, SAR_Rx: %h", w_SAR_Tx, w_SAR_Rx);
    else
      $display("Test Failed - Signatures Do Not Match. SAR_Tx: %h, SAR_Rx: %h", w_SAR_Tx, w_SAR_Rx);

    #1000;  // Add a delay to ensure the simulation runs long enough
    $finish();
  end

endmodule
*/

`timescale 1ns/1ps

module UART_TB;

  // Inputs
  reg clk;
  reg rst_n;
  reg mode;
  reg i_TX_DV;
  reg [7:0] tx_byte;
  reg [1:0] baud_rate;

  // Outputs
  wire o_RX_DV;
  wire [7:0] rx_byte;
  wire [15:0] o_SAR_Tx;
  wire [15:0] o_SAR_Rx;

  reg [4:0] i;

  // Instantiate the DUT (Device Under Test)
  UART_TOP uut (
    .clk(clk),
    .rst_n(rst_n),
    .mode(mode),
    .i_TX_DV(i_TX_DV),
    .tx_byte(tx_byte),
    .baud_rate(baud_rate),
    .o_RX_DV(o_RX_DV),
    .rx_byte(rx_byte),
    .o_SAR_Tx(o_SAR_Tx),
    .o_SAR_Rx(o_SAR_Rx)
  );

  // Clock generation: 50MHz
  always #10 clk = ~clk;

  // Task to send a byte
  task send_byte(input [7:0] data);
    begin
      tx_byte = data;
      i_TX_DV = 1;
      #20;
      i_TX_DV = 0;
    end
  endtask

  initial begin
    // Initialize inputs
    clk = 0;
    rst_n = 1;
    mode = 0;
    i_TX_DV = 0;
    tx_byte = 8'h00;
    baud_rate = 2'b10; // 9600 baud (adjusted for test)

    // Apply reset
    #100;
    rst_n = 0;
    // Wait for reset de-assertion
    #100;
    rst_n = 1;
    #10;

    // ------------ Manual Mode ------------
    //mode = 0;
    //$display("Manual Mode: Sending byte 0x55");
    //send_byte(8'h55);

    //wait (o_RX_DV == 1);
    //$display("Received Byte: %h | SAR_Tx: %d | SAR_Rx: %d", rx_byte, o_SAR_Tx, o_SAR_Rx);

    //#50000;

    // ------------ Test Mode (BIST) ------------
    mode = 1;
    for(i =0; i<10 ; i = i+1)
    begin
    $display("Test Mode (BIST): Sending LFSR-generated byte");
    send_byte(8'h00); // tx_byte ignored in test mode

    wait (o_RX_DV == 1);
    $display("Received Byte: %h | SAR_Tx: %d | SAR_Rx: %d", rx_byte, o_SAR_Tx, o_SAR_Rx);
    #5000;
    end
    //#50000;
    $display("Received Byte: %h | SAR_Tx: %d | SAR_Rx: %d", rx_byte, o_SAR_Tx, o_SAR_Rx);
    $display("Simulation completed.");
    $finish;
  end

  initial
  begin
    $dumpfile("dump.vcd");
    $dumpvars(0, UART_TB);
    //$dumpvars(1, UART_TX_INST);
    //$dumpvars(1, UART_RX_INST);
    end

endmodule
